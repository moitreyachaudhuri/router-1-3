module synchroniser(input clk,rstn,detect_add,write_enb_reg,full_0,full_1,full_2,read_enb_0,read_enb_1,read_enb_2,empty_0,empty_1,empty_2,input [1:0] data_in,output vld_out_0,vld_out_1,vld_out_2,output reg fifo_full,soft_reset_0,soft_reset_1,soft_reset_2,output reg [2:0] write_enb);
reg [1:0] int_add_reg;
reg timer_0,timer_1,timer_2;
always @(posedge clk)
begin
if (!rstn)
int_add_reg<=0;
else if(detect_add)
int_add_reg<=data_in;
end
//write_enable logic
always @(*)
begin
if (write_enb_reg)
	begin
	case(int_add_reg)
	2'b00: write_enb=3'b001;
	2'b01: write_enb=3'b010;
	2'b10: write_enb=3'b100;
	default: write_enb=3'b000;
	endcase
	end
end
//fifo_full logic
always @(*)
begin
	begin
	case(int_add_reg)
	2'b00: fifo_full=full_0;
	2'b01: fifo_full=full_1;
	2'b10: fifo_full=full_2;
	default: fifo_full=1'b0;
	endcase
	end
end
assign vld_out_0=~empty_0;
assign vld_out_1=~empty_1;
assign vld_out_2=~empty_2;
//timer_0 and soft_reset_0 logic
always @(posedge clk)
begin
	if (!rstn)
	begin
		timer_0<=0;
		soft_reset_0<=0;
	end
	else if(vld_out_0)
	begin
		if (!read_enb_0)
		begin
			if(timer_0==5'd29)
			begin
				soft_reset_0<=1'b1;
				timer_0<=0;
			end
			else	
			begin
				soft_reset_0<=0;
				timer_0<=timer_0+1'b1;
			end
		end
	end
end
always @(posedge clk)
begin
	if (!rstn)
	begin
		timer_1<=0;
		soft_reset_1<=0;
	end
	else if(vld_out_1)
	begin
		if (!read_enb_1)
		begin
			if(timer_1==5'd29)
			begin
				soft_reset_1<=1'b1;
				timer_1<=0;
			end
			else	
			begin
				soft_reset_1<=0;
				timer_1<=timer_1+1'b1;
			end
		end
	end
end
always @(posedge clk)
begin
	if (!rstn)
	begin
		timer_2<=0;
		soft_reset_2<=0;
	end
	else if(vld_out_2)
	begin
		if (!read_enb_2)
		begin
			if(timer_2==5'd29)
			begin
				soft_reset_2<=1'b1;
				timer_2<=0;
			end
			else	
			begin
				soft_reset_2<=0;
				timer_2<=timer_2+1'b1;
			end
		end
	end
end
	


endmodule